/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_APB_ENV_PKG_SVH
`define YUU_APB_ENV_PKG_SVH

  `include "yuu_apb_env_config.sv"
  `include "yuu_apb_env.sv"

`endif
