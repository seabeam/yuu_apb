/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_APB_COMMON_PKG_SVH
`define YUU_APB_COMMON_PKG_SVH

  `include "yuu_apb_type.sv"
  `include "yuu_apb_error.sv"
  `include "yuu_apb_item.sv"
  `include "yuu_apb_agent_config.sv"

`endif
