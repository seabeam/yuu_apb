/////////////////////////////////////////////////////////////////////////////////////
// Copyright 2019 seabeam@yahoo.com - Licensed under the Apache License, Version 2.0
// For more information, see LICENCE in the main folder
/////////////////////////////////////////////////////////////////////////////////////
`ifndef YUU_APB_COMMON_PKG
`define YUU_APB_COMMON_PKG

  `include "yuu_apb_type.svh"
  `include "yuu_apb_error.sv"
  `include "yuu_apb_item.sv"
  `include "yuu_apb_agent_config.sv"

`endif
